../../src/MOM6/ice_ocean_SIS2/OM4_025/INPUT/Faroe_GS_edits.cdl