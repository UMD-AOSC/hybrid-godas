../../../src/MOM6/ice_ocean_SIS2/OM4_025/INPUT/vgrid_75_2m_575m.cdl