../../../src/MOM6/ice_ocean_SIS2/OM4_025/INPUT/hycom1_75.cdl