../../../src/MOM6/ice_ocean_SIS2/OM4_025/INPUT/analysis_vgrid_lev35.v1.cdl